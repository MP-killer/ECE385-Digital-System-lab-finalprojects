module character_rom ( input [6:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
//left
16'b0000111111000000,
16'b0011111111110000,
16'b0111111111111000,
16'b0011111111111100,
16'b0001111111111110,
16'b0000111111111110,
16'b0000001111111110,
16'b0000000111111110,
16'b0000001111111110,
16'b0000111111111110,
16'b0001111111111110,
16'b0011111111111100,
16'b0111111111111000,
16'b0011111111110000,
16'b0001111111100000,
16'b0000111111000000,

//right
16'b0000001111110000,
16'b0000111111111100,
16'b0001111111111110,
16'b0011111111111100,
16'b0111111111111000,
16'b0111111111110000,
16'b0111111111000000,
16'b0111111110000000,
16'b0111111111000000,
16'b0111111111110000,
16'b0111111111111000,
16'b0011111111111100,
16'b0001111111111110,
16'b0000111111111100,
16'b0000011111111000,
16'b0000001111110000,
//down;
16'b0000000000000000,
16'b0000001111000000,
16'b0000111111110000,
16'b0011111111111100,
16'b0011111111111100,
16'b0111111111111110,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111001111111,
16'b1111111001111111,
16'b0111100000011110,
16'b0111000000001110,
16'b0010000000000100,
16'b0000000000000000,
16'b0000000000000000,
//up
16'b0000000000000000,
16'b0000000000000000,
16'b0010000000000100,
16'b0111000000001110,
16'b0111100000011110,
16'b1111111001111111,
16'b1111111001111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b0111111111111110,
16'b0011111111111100,
16'b0011111111111100,
16'b0000111111110000,
16'b0000001111000000,
16'b0000000000000000,

//ghost
16'b0000001111000000,
16'b0000111111110000,
16'b0011111111111100,
16'b0111111111111110,
16'b0111111111111110,
16'b0111111111111110,
16'b0111000110001110,
16'b1111000110001111,
16'b1111111111111111,
16'b1111111111111111,
16'b1000111000110001,
16'b1011000111001101,
16'b1111111111111111,
16'b1110111001110111,
16'b1100011001100011,
16'b1000001001000001,
        };

	assign data = ROM[addr];

endmodule  