module endscene_rom ( input [4:0]	addr,
						output[39:0] 	data
					 );
		parameter ADDR_WIDTH = 5;
   	parameter DATA_WIDTH =  40;			
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {

		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000011110000011100001100001101111111000,
		40'b0000110011000110110001110011100110011000,
		40'b0001100001001100011001111111100110001000,
		40'b0001100000001100011001111111100110100000,
		40'b0001100000001111111001101101100111100000,
		40'b0001101111001100011001101101100110100000,
		40'b0001100011001100011001100001100110000000,
		40'b0001100011001100011001100001100110001000,
		40'b0000110011001100011001100001100110011000,
		40'b0000011101001100011001100001101111111000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000111110001100001101111111001111110000,
		40'b0001100011001100001100110011000110011000,
		40'b0001100011001100001100110001000110011000,
		40'b0001100011001100001100110100000110011000,
		40'b0001100011001100001100111100000111110000,
		40'b0001100011001100001100110100000110110000,
		40'b0001100011001100001100110000000110011000,
		40'b0001100011000110011000110001000110011000,
		40'b0001100011000011110000110011000110011000,
		40'b0000111110000001100001111111001110011000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
		40'b0000000000000000000000000000000000000000,
 };

	assign data = ROM[addr];

endmodule






















