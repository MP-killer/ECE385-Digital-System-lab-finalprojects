module room_rom ( input [4:0]	addr,
						output[39:0] 	data
					 );
		parameter ADDR_WIDTH = 5;
   	parameter DATA_WIDTH =  40;			
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        40'b0000000000000000000000000000000000000000, // 0
		  40'b0000001111111111111111111111111111000000, // 1
        40'b0000001000000000000110000000000001000000, // 2
        40'b0000001011110111110110111110111101000000, // 3
        40'b0000001011110111110110111110111101000000, // 4
        40'b0000001000000000000000000000000001000000, // 5
        40'b0000001011110110111111110110111101000000, // 6
        40'b0000001000000110000110000110000001000000, // 7
        40'b0000001111110111110110111110111111000000, // 8
        40'b0000000000010111110110111110100000000000, // 9
		  40'b0000000000010110000000000110100000000000, // 10
		  40'b0000000000010110111111110110100000000000, // 11
        40'b0000001111110110100000010110111111000000, // 12
        40'b0000001000000000100000010000000001000000, // 13
        40'b0000001111110110100000010110111111000000, // 14
        40'b0000000000010110111111110110100000000000, // 15
        40'b0000000000010110000000000110100000000000, // 16
        40'b0000000000010110111111110110100000000000, // 17
        40'b0000001111110110111111110110111111000000, // 18
        40'b0000001000000000000110000000000001000000, // 19
		  40'b0000001011110111110110111110111101000000, // 20
		  40'b0000001000110000000000000000110001000000, // 21
        40'b0000001110110110111111110110110111000000, // 22
        40'b0000001110110110111111110110110111000000, // 23
        40'b0000001000000110000110000110000001000000, // 24
        40'b0000001011111111110110111111111101000000, // 25
        40'b0000001011111111110110111111111101000000, // 26
        40'b0000001000000000000000000000000001000000, // 27
        40'b0000001111111111111111111111111111000000, // 28
        40'b0000000000000000000000000000000000000000, // 29

        };

	assign data = ROM[addr];

endmodule

module room_rom_4 (  input [4:0]	addr1,
							input [4:0]	addr2,
							input [4:0]	addr3,
							input [4:0]	addr4,
						   output[39:0] 	data1,
						   output[39:0] 	data2,
						   output[39:0] 	data3,
						output[39:0] 	data4
					 );
		parameter ADDR_WIDTH = 5;
   	parameter DATA_WIDTH =  40;			
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        40'b0000000000000000000000000000000000000000, // 0
		  40'b0000001111111111111111111111111111000000, // 1
        40'b0000001000000000000110000000000001000000, // 2
        40'b0000001011110111110110111110111101000000, // 3
        40'b0000001011110111110110111110111101000000, // 4
        40'b0000001000000000000000000000000001000000, // 5
        40'b0000001011110110111111110110111101000000, // 6
        40'b0000001000000110000110000110000001000000, // 7
        40'b0000001111110111110110111110111111000000, // 8
        40'b0000000000010111110110111110100000000000, // 9
		  40'b0000000000010110000000000110100000000000, // 10
		  40'b0000000000010110111111110110100000000000, // 11
        40'b0000001111110110100000010110111111000000, // 12
        40'b0000001000000000100000010000000001000000, // 13
        40'b0000001111110110100000010110111111000000, // 14
        40'b0000000000010110111111110110100000000000, // 15
        40'b0000000000010110000000000110100000000000, // 16
        40'b0000000000010110111111110110100000000000, // 17
        40'b0000001111110110111111110110111111000000, // 18
        40'b0000001000000000000110000000000001000000, // 19
		  40'b0000001011110111110110111110111101000000, // 20
		  40'b0000001000110000000000000000110001000000, // 21
        40'b0000001110110110111111110110110111000000, // 22
        40'b0000001110110110111111110110110111000000, // 23
        40'b0000001000000110000110000110000001000000, // 24
        40'b0000001011111111110110111111111101000000, // 25
        40'b0000001011111111110110111111111101000000, // 26
        40'b0000001000000000000000000000000001000000, // 27
        40'b0000001111111111111111111111111111000000, // 28
        40'b0000000000000000000000000000000000000000, // 29

        };

	assign data1 = ROM[addr1];
	assign data2 = ROM[addr2];
	assign data3 = ROM[addr3];
	assign data4 = ROM[addr4];


endmodule

module room_rom_8 (  input [4:0]	addr1,
							input [4:0]	addr2,
							input [4:0]	addr3,
							input [4:0]	addr4,
							input [4:0]	addr5,
							input [4:0]	addr6,
							input [4:0]	addr7,
							input [4:0]	addr8,
						   output[39:0] 	data1,
						   output[39:0] 	data2,
						   output[39:0] 	data3,
						   output[39:0] 	data4,
							output[39:0] 	data5,
						   output[39:0] 	data6,
						   output[39:0] 	data7,
						   output[39:0] 	data8
					 );
		parameter ADDR_WIDTH = 5;
   	parameter DATA_WIDTH =  40;			
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        40'b0000000000000000000000000000000000000000, // 0
		  40'b0000001111111111111111111111111111000000, // 1
        40'b0000001000000000000110000000000001000000, // 2
        40'b0000001011110111110110111110111101000000, // 3
        40'b0000001011110111110110111110111101000000, // 4
        40'b0000001000000000000000000000000001000000, // 5
        40'b0000001011110110111111110110111101000000, // 6
        40'b0000001000000110000110000110000001000000, // 7
        40'b0000001111110111110110111110111111000000, // 8
        40'b0000000000010111110110111110100000000000, // 9
		  40'b0000000000010110000000000110100000000000, // 10
		  40'b0000000000010110111111110110100000000000, // 11
        40'b0000001111110110100000010110111111000000, // 12
        40'b0000001000000000100000010000000001000000, // 13
        40'b0000001111110110100000010110111111000000, // 14
        40'b0000000000010110111111110110100000000000, // 15
        40'b0000000000010110000000000110100000000000, // 16
        40'b0000000000010110111111110110100000000000, // 17
        40'b0000001111110110111111110110111111000000, // 18
        40'b0000001000000000000110000000000001000000, // 19
		  40'b0000001011110111110110111110111101000000, // 20
		  40'b0000001000110000000000000000110001000000, // 21
        40'b0000001110110110111111110110110111000000, // 22
        40'b0000001110110110111111110110110111000000, // 23
        40'b0000001000000110000110000110000001000000, // 24
        40'b0000001011111111110110111111111101000000, // 25
        40'b0000001011111111110110111111111101000000, // 26
        40'b0000001000000000000000000000000001000000, // 27
        40'b0000001111111111111111111111111111000000, // 28
        40'b0000000000000000000000000000000000000000, // 29

        };

	assign data1 = ROM[addr1];
	assign data2 = ROM[addr2];
	assign data3 = ROM[addr3];
	assign data4 = ROM[addr4];
	assign data5 = ROM[addr5];
	assign data6 = ROM[addr6];
	assign data7 = ROM[addr7];
	assign data8 = ROM[addr8];

endmodule


module room_rom_10 ( input [4:0]	addr1,
							input [4:0]	addr2,
							input [4:0]	addr3,
							input [4:0]	addr4,
							input [4:0]	addr5,
							input [4:0]	addr6,
							input [4:0]	addr7,
							input [4:0]	addr8,
							input [4:0] addr9,
							input [4:0] addr10,
						   output[39:0] 	data1,
						   output[39:0] 	data2,
						   output[39:0] 	data3,
						   output[39:0] 	data4,
							output[39:0] 	data5,
						   output[39:0] 	data6,
						   output[39:0] 	data7,
						   output[39:0] 	data8,
						   output[39:0] 	data9,
						   output[39:0] 	data10
					 );
		parameter ADDR_WIDTH = 5;
   	parameter DATA_WIDTH =  40;			
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        40'b0000000000000000000000000000000000000000, // 0
		  40'b0000001111111111111111111111111111000000, // 1
        40'b0000001000000000000110000000000001000000, // 2
        40'b0000001011110111110110111110111101000000, // 3
        40'b0000001011110111110110111110111101000000, // 4
        40'b0000001000000000000000000000000001000000, // 5
        40'b0000001011110110111111110110111101000000, // 6
        40'b0000001000000110000110000110000001000000, // 7
        40'b0000001111110111110110111110111111000000, // 8
        40'b0000000000010111110110111110100000000000, // 9
		  40'b0000000000010110000000000110100000000000, // 10
		  40'b0000000000010110111111110110100000000000, // 11
        40'b0000001111110110100000010110111111000000, // 12
        40'b0000001000000000100000010000000001000000, // 13
        40'b0000001111110110100000010110111111000000, // 14
        40'b0000000000010110111111110110100000000000, // 15
        40'b0000000000010110000000000110100000000000, // 16
        40'b0000000000010110111111110110100000000000, // 17
        40'b0000001111110110111111110110111111000000, // 18
        40'b0000001000000000000110000000000001000000, // 19
		  40'b0000001011110111110110111110111101000000, // 20
		  40'b0000001000110000000000000000110001000000, // 21
        40'b0000001110110110111111110110110111000000, // 22
        40'b0000001110110110111111110110110111000000, // 23
        40'b0000001000000110000110000110000001000000, // 24
        40'b0000001011111111110110111111111101000000, // 25
        40'b0000001011111111110110111111111101000000, // 26
        40'b0000001000000000000000000000000001000000, // 27
        40'b0000001111111111111111111111111111000000, // 28
        40'b0000000000000000000000000000000000000000, // 29

        };

	assign data1 = ROM[addr1];
	assign data2 = ROM[addr2];
	assign data3 = ROM[addr3];
	assign data4 = ROM[addr4];
	assign data5 = ROM[addr5];
	assign data6 = ROM[addr6];
	assign data7 = ROM[addr7];
	assign data8 = ROM[addr8];
	assign data9 = ROM[addr9];
	assign data10 = ROM[addr10];

endmodule
